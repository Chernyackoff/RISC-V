LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Adder IS
    GENERIC (ADDER_DATA_WIDTH : INTEGER := 32);
    PORT (
        ADDER_INPUT_A : IN UNSIGNED(ADDER_DATA_WIDTH - 1 DOWNTO 0);
        ADDER_INPUT_B : IN UNSIGNED(ADDER_DATA_WIDTH - 1 DOWNTO 0);
        ADDER_OUTPUT : OUT UNSIGNED(ADDER_DATA_WIDTH - 1 DOWNTO 0)
    );
END ENTITY Adder;

ARCHITECTURE RTL OF Adder IS
BEGIN
    ADDER_OUTPUT <= ADDER_INPUT_A + ADDER_INPUT_B;
END ARCHITECTURE RTL;